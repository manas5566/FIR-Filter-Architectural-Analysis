module Carryskip_32(s, Cout, x, y, Cin);
  input [31:0] x, y;
  output [31:0] s;
  output Cout;
  input Cin;
  wire [31:0] C, p;
  wire pout;
  fa f1(x[0], y[0], Cin, s[0], C[0], p[0]);
  fa f2(x[1], y[1], C[0], s[1], C[1], p[1]);
  fa f3(x[2], y[2], C[1], s[2], C[2], p[2]);
  fa f4(x[3], y[3], C[2], s[3], C[3], p[3]);
  fa f5(x[4], y[4], C[3], s[4], C[4], p[4]);
  fa f6(x[5], y[5], C[4], s[5], C[5], p[5]);
  fa f7(x[6], y[6], C[5], s[6], C[6], p[6]);
  fa f8(x[7], y[7], C[6], s[7], C[7], p[7]);
  fa f9(x[8], y[8], C[7], s[8], C[8], p[8]);
  fa f10(x[9], y[9], C[8], s[9], C[9], p[9]);
  fa f11(x[10], y[10], C[9], s[10], C[10], p[10]);
  fa f12(x[11], y[11], C[10], s[11], C[11], p[11]);
  fa f13(x[12], y[12], C[11], s[12], C[12], p[12]);
  fa f14(x[13], y[13], C[12], s[13], C[13], p[13]);
  fa f15(x[14], y[14], C[13], s[14], C[14], p[14]);                           
  fa f16(x[15], y[15], C[14], s[15], C[15], p[15]);
  fa f17(x[16], y[16], C[15], s[16], C[16], p[16]);
  fa f18(x[17], y[17], C[16], s[17], C[17], p[17]);
  fa f19(x[18], y[18], C[17], s[18], C[18], p[18]);
  fa f20(x[19], y[19], C[18], s[19], C[19], p[19]);
  fa f21(x[20], y[20], C[19], s[20], C[20], p[20]);
  fa f22(x[21], y[21], C[20], s[21], C[21], p[21]);
  fa f23(x[22], y[22], C[21], s[22], C[22], p[22]);
  fa f24(x[23], y[23], C[22], s[23], C[23], p[23]);
  fa f25(x[24], y[24], C[23], s[24], C[24], p[24]);
  fa f26(x[25], y[25], C[24], s[25], C[25], p[25]);
  fa f27(x[26], y[26], C[25], s[26], C[26], p[26]);
  fa f28(x[27], y[27], C[26], s[27], C[27], p[27]);
  fa f29(x[28], y[28], C[27], s[28], C[28], p[28]);
  fa f30(x[29], y[29], C[28], s[29], C[29], p[29]);
  fa f31(x[30], y[30], C[29], s[30], C[30], p[30]);
  fa f32(x[31], y[31], C[30], s[31], C[31], p[31]);
  assign pout= ( p[0]& p[1] & p[2] & p[3] & p[4]& p[5] & p[6] & p[7] & p[8]& p[9] & p[10]& p[11] & p[12] & p[13] & p[14]& p[15] & p[16] & p[17] & p[18]& p[19] & p[20]& p[21] & p[22] & p[23] & p[24]& p[25] & p[26] & p[27] & p[28]& p[29] & p[30] & p[31]);
  mux2_1 m1(C[31], Cin, pout , Cout);
endmodule